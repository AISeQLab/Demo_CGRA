`define LDM_DEPTH 24
`define CTX_RC_DEPTH 1072
`define CTX_PE_DEPTH 1072
`define CTX_IM_DEPTH 1072
